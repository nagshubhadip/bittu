module muxtb;
reg s;
reg [3:0]d1;
reg [3:0]d0;
wire [3:0]f;
mux4bit m1(f,s,d1,d0);
initial
	begin
	s=0;d1=4'bxxxx;d0=4'b0000;
	#5 d0=4'b0001;
	#5 d0=4'b0010;
	#5 d0=4'b0011;
	#5 d0=4'b0100;
	#5 d0=4'b0101;
	#5 d0=4'b0110;
	#5 d0=4'b0111;
	#5 d0=4'b1000;
	#5 d0=4'b1001;
	#5 d0=4'b1010;
	#5 d0=4'b1011;
	#5 d0=4'b1100;
	#5 d0=4'b1101;
	#5 d0=4'b1110;
	#5 d0=4'b1111;
	#5 s=1;d1=4'b0000;d0=4'bxxxx;
	#5 d1=4'b0001;
	#5 d1=4'b0010;
	#5 d1=4'b0011;
	#5 d1=4'b0100;
	#5 d1=4'b0101;
	#5 d1=4'b0110;
	#5 d1=4'b0111;
	#5 d1=4'b1000;
	#5 d1=4'b1001;
	#5 d1=4'b1010;
	#5 d1=4'b1011;
	#5 d1=4'b1100;
	#5 d1=4'b1101;
	#5 d1=4'b1110;
	#5 d1=4'b1111;
	end
initial 
	begin
	$monitor (" s = %b   D1 = %b  D0 = %b   F = %b ",s,d1,d0,f);
	end
endmodule
